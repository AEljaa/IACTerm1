module top #(
    parameter D_WIDTH=8,
              C_WIDTH=16
)(
input logic clk, //clk
input logic trigger,//trigger
input logic rst, //reset
input  logic [C_WIDTH-1:0] N,     	 // clock divided by N+1
output logic [D_WIDTH-1:0] data_out //semi random output
);


logic tick_time; //interconnect gerated tick wire from the clktick module output

logic cmd_seq; //result from our f1_fsm of wheter we use the clock tick or delay signal (if 1 then use)

logic cmd_delay; //the value we feed into the trigger value in our delay module

logic random_num;//random num from our lfsr_7b modle that we cary over to our delay module

logic time_out;// the delayed time out signal we feed into the 0 of our mux

logic mux_val;


assign mux_val = cmd_seq ? tick_time : time_out ;

f1_fsm  f1_lights (
    .clk (clk),
    .en  (mux_val),
    .rst (rst),
    .trigger(trigger),
    .cmd_seq(cmd_seq),//output fed into mux as selector and the en of clktick
    .cmd_delay(cmd_delay),//output we feed into the trigger value of delay module
    .data_out (data_out)//output the sequnce we see
);


clktick clocktick(
    .clk (clk),
    .N   (N),
    .en (cmd_seq),
    .rst (rst),
    .tick (tick_time)//output we feed into mux
);

lfsr_7b lfsr (
    .clk(clk),
    .rst(rst),
    .data_out(random_num)//output psuedo random number generated by our lfsr
);

delay delay(
    .clk(clk),
    .rst(rst),
    .trigger(cmd_delay),
    .n(random_num),
    .time_out(time_out)
);

endmodule

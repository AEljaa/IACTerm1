module counter_flg #(
    parameter WIDTH = 8 
)

(
    //Interface Signals
    input logic clk, //clock
    input logic rst, //reset
    input logic en, //enable
    output logic [WIDTH-1:0] count //count output
);

always_ff @(posedge clk) 
    if (rst) count <= {WIDTH{1'b0}}; 
    else if (en)  count <= count + {{WIDTH-1{1'b0}},1'b1};
    else count <= count - {{WIDTH-1{1'b0}},1'b1};

endmodule;
 

module top #(
    parameter D_WIDTH=8,
              C_WIDTH=16
)(
input logic clk, //clk
input logic trigger,//trigger
input logic rst, //reset
input  logic [C_WIDTH-1:0] N,     	 // clock divided by N+1
output logic [D_WIDTH-1:0] data_out //semi random output
);


logic tick_time; //interconnect gerated tick wire from the clktick module output

logic cmd_seq=1'b1; //result from our f1_fsm of wheter we use the clock tick or delay signal (if 1 then use/1 by default)

logic cmd_delay=1'b0; //the value we feed into the trigger value in our delay module (0 by default)

logic [6:0] random_num;//random num from our lfsr_7b modle that we cary over to our delay module

logic delay_time;// the delayed time out signal we feed into the 0 of our mux




f1_fsm  f1_lights (
    .clk (clk),
    .en  (cmd_seq ? tick_time : delay_time),
    .rst (rst),
    .trigger(trigger),
    .cmd_seq(cmd_seq),//output fed into mux as selector and the en of clktick
    .cmd_delay(cmd_delay),//output we feed into the trigger value of delay module
    .data_out (data_out)//output the sequnce we see
);


clktick clocktick(
    .clk (clk),
    .N   (N),
    .en (cmd_seq),
    .rst (rst),
    .tick (tick_time)//output we feed into mux
);

lfsr_7b lfsr(
    .clk(clk),
    .rst(rst),
    .data_out(random_num)//output psuedo random number generated by our lfsr
);

delay delay(
    .clk(clk),
    .rst(rst),
    .trigger(cmd_delay),
    .n(random_num),
    .time_out(delay_time)
);

endmodule

module lfsr_7b (
    input logic clk,
    input logic rst,
    output logic [7:1] data_out //semi random output
);

logic [7:1] sreg;

always_ff @(posedge clk, posedge rst) begin
    if (rst)
        sreg <= 7'b1;
    else 
        sreg <= {sreg[6:1], sreg[7] ^ sreg[3]};

    assign data_out = sreg ;
end
endmodule

